library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity NIVEL is
    Port ( CLK : in  STD_LOGIC;
           CLR : in  STD_LOGIC;
           NIV_ALTO : out  STD_LOGIC);
end NIVEL;

architecture DETECTOR of NIVEL is
SIGNAL PCLK, NCLK: STD_LOGIC;
begin

	PPCLK: PROCESS(CLK,CLR)
	BEGIN
		IF(CLR = '1') THEN
			PCLK<='0';
		ELSIF(RISING_EDGE(CLK))THEN
			PCLK<=NOT PCLK;
		END IF;
	END PROCESS PPCLK;
	
	NIV_ALTO<=PCLK XOR NCLK;
	
	PNCLK: PROCESS(CLK,CLR)
	BEGIN
		IF(CLR = '1') THEN
			NCLK<='0';
		ELSIF(FALLING_EDGE(CLK))THEN
			NCLK<=NOT NCLK;
		END IF;
	END PROCESS PNCLK;

end DETECTOR;

