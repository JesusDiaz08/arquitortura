library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FUNCION is
    Port ( A : in  STD_LOGIC_VECTOR (3 downto 0);
           D : out STD_LOGIC_VECTOR (19 downto 0));
end FUNCION;

architecture MEMORIA of FUNCION is

	TYPE ROM IS ARRAY (0 TO 2**4) OF STD_LOGIC_VECTOR(D' RANGE);
	
	CONSTANT MEM_FUN : ROM := (
		--12345678901234567890
		"00000100110000011001",	--ADD
		"00000100110000111001",	--SUB
		"00000100110000000001",	--AND
		"00000100110000001001",	--OR
		"00000100110000010001",	--XOR
		"00000100110001101001",	--NAND
		"00000100110001100001",	--NOR
		"00000100110000110001",	--XNOR
		"00000100110001101001",	--NOT
		"00000011100000000000",	--SLL 
		"00000010100000000000",	--SRL 
		OTHERS => (OTHERS => '0')		
	);

begin
	D 	<=	MEM_FUN(0) WHEN 	A="0000" ELSE
			MEM_FUN(1) WHEN 	A="0001" ELSE
			MEM_FUN(2) WHEN 	A="0010" ELSE
			MEM_FUN(3) WHEN 	A="0011" ELSE
			MEM_FUN(4) WHEN 	A="0100" ELSE
			MEM_FUN(5) WHEN 	A="0101" ELSE
			MEM_FUN(6) WHEN 	A="0110" ELSE
			MEM_FUN(7) WHEN 	A="0111" ELSE
			MEM_FUN(8) WHEN 	A="1000" ELSE
			MEM_FUN(9) WHEN 	A="1001" ELSE
			MEM_FUN(10) WHEN 	A="1010" ELSE
			MEM_FUN(11) WHEN 	A="1011" ELSE
			MEM_FUN(12);
end MEMORIA;