library IEEE;
library WORK;
use IEEE.STD_LOGIC_1164.all;
use WORK.MI_PAQUETE.all;

entity main is
    Port ( DATOS : in  STD_LOGIC_VECTOR (7 downto 0);
           INI : in  STD_LOGIC;
           CLR : in  STD_LOGIC;
           CLK : in  STD_LOGIC;
           DISP : out  STD_LOGIC_VECTOR (6 downto 0));
end main;

architecture Behavioral of main is
--CONSTANTES
CONSTANT DIG0 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
CONSTANT DIG1 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
CONSTANT DIG2 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
CONSTANT DIG3 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
CONSTANT DIG4 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001100";
CONSTANT DIG5 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
CONSTANT DIG6 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100000";
CONSTANT DIG7 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001110";
CONSTANT DIG8 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
CONSTANT DIG9 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001100";
CONSTANT DIGA : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001000";
CONSTANT DIGB : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1100000";
CONSTANT DIGC : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000";
CONSTANT DIGD : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1000010";
CONSTANT DIGE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000";
CONSTANT DIGF : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0111000";
--SE�ALES
signal QB, E:STD_LOGIC_VECTOR(3 DOWNTO 0);
signal QA:STD_LOGIC_VECTOR(7 DOWNTO 0);
signal LB, IB, LA, EA, SD, Z: STD_LOGIC;
--signal SAL: STD_LOGIC_VECTOR(6 DOWNTO 0);


begin
	CONT: contador PORT MAP(X"0", QB, LB, IB, CLK, CLR);
	REG: registro PORT MAP(DATOS, QA, LA, EA, CLK, CLR);
	COD: codigo PORT MAP(E, DISP); --NOSE CUAL SEA LA SALIDA
	CON: control PORT MAP(CLK, CLR, INI, Z, QA(0), LA, SH, LB, IB, SD);--CHECAR QUIEN ES A0

	--DISP<=DIG0 WHEN (SD = '0') ELSE
	--		DIG1 WHEN (QA = '1');
	

	--COMPUERTA DE BANDERA Z
end Behavioral;

