--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package mi_paquete is

-- type <new_type> is
--  record
--    <type_name>        : std_logic_vector( 7 downto 0);
--    <type_name>        : std_logic;
-- end record;
--
-- Declare constants
--
-- constant <constant_name>		: time := <time_unit> ns;
-- constant <constant_name>		: integer := <value;
--
-- Declare functions and procedure
--
-- function <function_name>  (signal <signal_name> : in <type_declaration>) return <type_declaration>;
-- procedure <procedure_name> (<type_declaration> <constant_name>	: in <type_declaration>);
--

end mi_paquete;

package body mi_paquete is

--component contador is
--    Port ( D : in  STD_LOGIC_VECTOR (3 downto 0);
--           Q : inout  STD_LOGIC_VECTOR (3 downto 0);
--           L : in  STD_LOGIC;
--           I : in  STD_LOGIC;
--           CLK : in  STD_LOGIC;
--           CLR : in  STD_LOGIC);
--end component;
 
end mi_paquete;
